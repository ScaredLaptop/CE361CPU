module IExecute(
    
    input clk,
    input rst,
);
endmodule // IExecute